
module fpga_rs232 (
	
	input  clk,
	input  rst_n,
	
	input  uart_rxd,
	output uart_txd
	);

	
	
	
	
endmodule	
