library verilog;
use verilog.vl_types.all;
entity tb_hsc is
end tb_hsc;
